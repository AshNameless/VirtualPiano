---------------------------------------------------------------------------------
---------------------------------------------------------------------------------
--predictor
--
-- 功能: 从二值化模块获取输入像素信息, 产生24位按键信号.
--
-- 描述: 第一个版本进行简单的监测, 检测到两个连续的1之后便计算当前像素的坐标, 并将对应的
--       按键位置位.
---------------------------------------------------------------------------------
---------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.constants.all;
-------------------------------------------------------
-------------------------------------------------------
entity predictor is 
generic(
	key_num : integer := 24;
);
port(
	rst_n : in std_logic;
	
	--输入像素信息. 由于经过二值化处理, 只有一位
	pixel : in std_logic;
	fsyn : in std_logic;  --帧同步
	pclk : in std_logic;  --像素时钟
	
	--输出按键信息
	key_statuses : out std_logic_vector()
	
	
);
end entity predictor;
-------------------------------------------------------
-------------------------------------------------------




