-------------------------------------------------------------------------
-------------------------------------------------------------------------
--fifo2sdram
--
-- 功能: 将fifo数据保存到sdram中
--
-- 描述: 只保留24位信息中最高位的1, 只保留一个音符. 再将转换后的单音符信息
--       作为选择器的输入, 选择对应的NCO相位步长, 并将其输出. 同时产生note_on
--       note_change等信号. 通过对比当前音符和上一音符来判断note_change是否该
--       置位, 由当前音符是否变为0来判断是否松键.
-------------------------------------------------------------------------
-------------------------------------------------------------------------